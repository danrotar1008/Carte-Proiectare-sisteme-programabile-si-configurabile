��- - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
 - -   C o m p a n y :    
 - -   E n g i n e e r :    
 - -    
 - -   C r e a t e   D a t e :         0 9 : 4 7 : 0 9   1 0 / 1 4 / 2 0 2 1    
 - -   D e s i g n   N a m e :    
 - -   M o d u l e   N a m e :         f s m 1   -   B e h a v i o r a l    
 - -   P r o j e c t   N a m e :    
 - -   T a r g e t   D e v i c e s :    
 - -   T o o l   v e r s i o n s :    
 - -   D e s c r i p t i o n :    
 - -  
 - -   D e p e n d e n c i e s :    
 - -  
 - -   R e v i s i o n :    
 - -   R e v i s i o n   0 . 0 1   -   F i l e   C r e a t e d  
 - -   A d d i t i o n a l   C o m m e n t s :    
 - -  
 - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
 l i b r a r y   I E E E ;  
 u s e   I E E E . S T D _ L O G I C _ 1 1 6 4 . A L L ;  
  
 - -   U n c o m m e n t   t h e   f o l l o w i n g   l i b r a r y   d e c l a r a t i o n   i f   u s i n g  
 - -   a r i t h m e t i c   f u n c t i o n s   w i t h   S i g n e d   o r   U n s i g n e d   v a l u e s  
 - - u s e   I E E E . N U M E R I C _ S T D . A L L ;  
  
 - -   U n c o m m e n t   t h e   f o l l o w i n g   l i b r a r y   d e c l a r a t i o n   i f   i n s t a n t i a t i n g  
 - -   a n y   X i l i n x   p r i m i t i v e s   i n   t h i s   c o d e .  
 - - l i b r a r y   U N I S I M ;  
 - - u s e   U N I S I M . V C o m p o n e n t s . a l l ;  
  
 e n t i t y   f s m 1   i s  
         P o r t   (   c l k   :   i n     S T D _ L O G I C ;  
                       r e s e t   :   i n     S T D _ L O G I C ;  
                       s w   :   i n     S T D _ L O G I C _ V E C T O R   ( 7   d o w n t o   0 ) ;  
                       l e d   :   o u t     S T D _ L O G I C _ V E C T O R   ( 7   d o w n t o   0 ) ) ;  
 e n d   f s m 1 ;  
  
 a r c h i t e c t u r e   B e h a v i o r a l   o f   f s m 1   i s  
  
       - - U t i l i z a i   n u m e   d e s c r i p t i v e   p e n t r u   s t r i ,   c u m   a r   f i   s t 1 _ r e s e t ,   s t 2 _ s e a r c h  
         t y p e   s t a t e _ t y p e   i s   ( s t 1 _ s t a r t ,   s t 2 _ 1 ,   s t 3 _ 2 ,   s t 4 _ 3 ) ;    
         s i g n a l   s t a t e ,   n e x t _ s t a t e   :   s t a t e _ t y p e ;      
       - - D e c l a r a i   s e m n a l e   i n t e r n e   p e n t r u   t o a t e   i e i r i l e   m a i n i i   d e   s t a r e  
 	   s i g n a l   l e d _ i   :   s t d _ l o g i c _ v e c t o r ( 7   d o w n t o   0 ) ;  
       - - a l t e   i e i r i  
  
 b e g i n  
  
       S Y N C _ P R O C :   p r o c e s s   ( c l k )  
       b e g i n  
             i f   ( c l k ' e v e n t   a n d   c l k   =   ' 1 ' )   t h e n  
                   i f   ( r e s e t   =   ' 1 ' )   t h e n  
                         s t a t e   < =   s t 1 _ s t a r t ;  
                         l e d   < =   " 0 0 0 0 0 0 0 0 " ;  
                   e l s e  
                         s t a t e   < =   n e x t _ s t a t e ;  
                         l e d   < =   l e d _ i ;  
                   e n d   i f ;                  
             e n d   i f ;  
       e n d   p r o c e s s ;  
    
       - - M a i n a   c u   s t r i   M O O R E   -   I e i r i   b a z a t e   n u m a i   p e   s t a r e  
       O U T P U T _ D E C O D E :   p r o c e s s   ( s t a t e )  
       b e g i n  
             - - i n t r o d u c e i   i n s t r u c i u n i   p e n t r u   a   d e c o d a   s e m n a l e l e   d e   i e i r e   i n t e r n e  
             i f   s t a t e   =   s t 1 _ s t a r t   t h e n  
                   l e d _ i   < =   " 1 0 0 0 0 0 0 1 " ;  
             e n d   i f ;  
             i f   s t a t e   =   s t 2 _ 1   t h e n  
                   l e d _ i   < =   " 1 1 1 1 0 0 0 0 " ;  
             e n d   i f ;  
             i f   s t a t e   =   s t 3 _ 2   t h e n  
                   l e d _ i   < =   " 1 1 0 0 1 1 0 0 " ;  
             e n d   i f ;  
             i f   s t a t e   =   s t 4 _ 3   t h e n  
                   l e d _ i   < =   " 1 0 1 0 1 0 1 0 " ;  
             e n d   i f ;  
       e n d   p r o c e s s ;  
    
       N E X T _ S T A T E _ D E C O D E :   p r o c e s s   ( s t a t e ,   s w )  
       b e g i n  
             - - d e c l a r a i   s t a r e a   i m p l i c i t   p e n t r u   n e x t _ s t a t e   p e n t r u   a   e v i t a   b l o c r i l e    
 	 	 n e x t _ s t a t e   < =   s t a t e ;   - - i m p l i c i t   e s t e   s   r m � i   � n   s t a r e a   a c t u a l  
             - - i n s e r e a z   i n s t r u c i u n i   p e n t r u   a   d e c o d a   n e x t _ s t a t e  
             c a s e   ( s t a t e )   i s  
                   w h e n   s t 1 _ s t a r t   = >  
                         i f   s w   =   " 0 0 0 0 0 0 0 1 "   t h e n  
                               n e x t _ s t a t e   < =   s t 2 _ 1 ;  
 	 	 	 	 e l s e  
 	 	 	 	 	 n e x t _ s t a t e   < =   s t 1 _ s t a r t ;  
                         e n d   i f ;  
                   w h e n   s t 2 _ 1   = >  
                         i f   s w   =   " 0 0 0 0 0 0 1 0 "   t h e n  
                               n e x t _ s t a t e   < =   s t 3 _ 2 ;  
 	 	 	 	 e l s i f   s w   =   " 0 0 0 0 0 0 1 1 "   t h e n  
 	 	 	 	 	 n e x t _ s t a t e   < =   s t 4 _ 3 ;  
 	 	 	 	 e l s e  
 	 	 	 	 	 n e x t _ s t a t e   < =   s t 2 _ 1 ;  
                         e n d   i f ;  
                   w h e n   s t 3 _ 2   = >  
 	 	 	 	 i f   s w   =   " 0 0 0 0 0 1 0 0 "   t h e n  
 	 	 	 	 	 n e x t _ s t a t e   < =   s t 1 _ s t a r t ;  
 	 	 	 	 e l s e  
 	 	 	 	 	 n e x t _ s t a t e   < =   s t 3 _ 2 ;  
 	 	 	 	 e n d   i f ;  
                   w h e n   s t 4 _ 3   = >  
 	 	 	 	 i f   s w   =   " 0 0 0 0 0 1 0 0 "   t h e n  
 	 	 	 	 	 n e x t _ s t a t e   < =   s t 1 _ s t a r t ;  
 	 	 	 	 e l s e  
 	 	 	 	 	 n e x t _ s t a t e   < =   s t 4 _ 3 ;  
 	 	 	 	 e n d   i f ;  
                   w h e n   o t h e r s   = >  
                         n e x t _ s t a t e   < =   s t 1 _ s t a r t ;  
             e n d   c a s e ;              
       e n d   p r o c e s s ;  
  
 e n d   B e h a v i o r a l ;  
  
 